module hole_number (
	input logic clk,
	input logic [10:0] pixelX,
	input logic [10:0] pixelY,
	input logic [2:0] holeNumber,
	output logic drawingRequestHoleNumber,
	output logic [7:0] RGBHoleNumber
);

const logic [7:0] TRANSPARENT_ENCODING = 8'hFF;
parameter int TOP_OFFSET = 0, DOWN_OFFSET = 479, LEFT_OFFSET = 0, RIGHT_OFFSET = 639;

// Because we use here a 32x16 bitmap and not 32x32 bitmap, we need to add an offset in order to center the number inside the hole
const int BITMAP_HEIGHT = 32;
const int BITMAP_WIDTH = 16;

const logic [10:0] LEFT_PLACE = LEFT_OFFSET - BITMAP_WIDTH / 2;
const logic [10:0] MIDDLE_PLACE = (LEFT_OFFSET + RIGHT_OFFSET) / 2 - BITMAP_WIDTH / 2;
const logic [10:0] RIGHT_PLACE = RIGHT_OFFSET - BITMAP_WIDTH / 2;
const logic [10:0] TOP_PLACE = TOP_OFFSET - BITMAP_HEIGHT / 2;
const logic [10:0] DOWN_PLACE = DOWN_OFFSET - BITMAP_HEIGHT / 2;

logic [10:0] holeTopLeftX, holeTopLeftY;

bit [0:5] [0:31] [0:15] NUMBER_BITMAP = {																	
{16'b	0000000011100000,
16'b	0000000111100000,
16'b	0000011111100000,
16'b	0000111111100000,
16'b	0001111111100000,
16'b	0011111111100000,
16'b	0111111011100000,
16'b	0111100011100000,
16'b	0111000011100000,
16'b	0010000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111},
									
{16'b	0000111111100000,
16'b	0001111111110000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000011111100,
16'b	1110000001111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000001111100,
16'b	0000000001111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011110000,
16'b	0000000011100000,
16'b	0000000111000000,
16'b	0000001111000000,
16'b	0000011110000000,
16'b	0000111100000000,
16'b	0001111100000000,
16'b	0001111100000000,
16'b	0011111000000000,
16'b	0111110000000001,
16'b	1111100000000011,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111},
																	
{16'b	0000111111100000,
16'b	0001111111111000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000001111100,
16'b	1110000001111100,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0001111111110000,
16'b	0001111111000000,
16'b	0001111111111000,
16'b	0001111111111000,
16'b	0000000011111100,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000111111,
16'b	1110000001111110,
16'b	1111100011111110,
16'b	1111111111111100,
16'b	1111111111111000,
16'b	0111111111111000,
16'b	0001111111000000},
																	
{16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000111111000,
16'b	0000001111111000,
16'b	0000001101111000,
16'b	0000011101111000,
16'b	0000011101111000,
16'b	0000111101111000,
16'b	0001111101111000,
16'b	0001111101111000,
16'b	0001111001111000,
16'b	0011111001111000,
16'b	0011110001111000,
16'b	0111100001111000,
16'b	0111100001111000,
16'b	1111000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000011111100},
																	
{16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111110,
16'b	0111111111111100,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111111111100000,
16'b	0111111111111000,
16'b	0111111111111000,
16'b	0111111111111100,
16'b	0010000011111110,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	1000000000111110,
16'b	1100000001111110,
16'b	1111100011111100,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	0001111111000000},
																	
{16'b	0000000111111100,
16'b	0000011111111110,
16'b	0000111111111110,
16'b	0001111111111111,
16'b	0001111100001111,
16'b	0011111100000001,
16'b	0011111000000000,
16'b	0111110000000000,
16'b	0111100000000000,
16'b	1111100000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111001111111000,
16'b	1111111111111100,
16'b	1111111111111110,
16'b	1111111111111111,
16'b	1111111101111111,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111100000001111,
16'b	1111100000001111,
16'b	0111110000011111,
16'b	0111111101111110,
16'b	0011111111111110,
16'b	0001111111111100,
16'b	0001111111111000,
16'b	0000011111100000}}; 


always_ff @(posedge clk)
begin 
	drawingRequestHoleNumber <= 1'b0;

	case(holeNumber)
		1: begin
			holeTopLeftX <= LEFT_PLACE;
			holeTopLeftY <= TOP_PLACE;	
			end		
		2: begin
			holeTopLeftX <= MIDDLE_PLACE;
			holeTopLeftY <= TOP_PLACE;	
			end
		3: begin
			holeTopLeftX <= RIGHT_PLACE;
			holeTopLeftY <= TOP_PLACE;	
			end
		4: begin
			holeTopLeftX <= RIGHT_PLACE;
			holeTopLeftY <= DOWN_PLACE;	
			end
		5: begin
			holeTopLeftX <= MIDDLE_PLACE;
			holeTopLeftY <= DOWN_PLACE;	
		end
		6: begin
			holeTopLeftX <= LEFT_PLACE;
			holeTopLeftY <= DOWN_PLACE;	
		end
	endcase

	if ((holeTopLeftX <= pixelX) && (holeTopLeftX + BITMAP_WIDTH > pixelX) && (holeTopLeftY + BITMAP_HEIGHT > pixelY) && (holeTopLeftY <= pixelY)) begin 
		drawingRequestHoleNumber <= NUMBER_BITMAP[holeNumber - 1][pixelY - holeTopLeftY][pixelX - holeTopLeftX];
	end
end  

assign RGBHoleNumber = TRANSPARENT_ENCODING - drawingRequestHoleNumber;

endmodule
