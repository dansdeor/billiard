module hole_collision (
					input logic clk,
					input logic resetN
);


endmodule
