module ball_draw (					
					output logic drawingRequestBall,
					output logic [7:0] RGBoutBall
);


endmodule
