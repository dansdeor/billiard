module statistics(
	input logic clk,
	
	input logic [10:0] pixelX,
	input logic [10:0] pixelY,
	
	input logic [7:0] score,
	input logic [7:0] attempts,
	
	input gameFinished,
	
	output logic drawingRequestStat,
	output logic [7:0] RGBoutStat
);

parameter int TOP_OFFSET = 0, DOWN_OFFSET = 479, LEFT_OFFSET = 0, RIGHT_OFFSET = 639;

const logic [10:0] MIDDLE_OFFSET_Y = (TOP_OFFSET + DOWN_OFFSET) / 2;
const logic [10:0] ATTEMPTS_OFFSET_X = (LEFT_OFFSET + RIGHT_OFFSET) / 8;
const logic [10:0] SCORE_OFFSET_X = 5 * (LEFT_OFFSET + RIGHT_OFFSET) / 8;

const int DIGIT_HEIGHT = 32;
const int DIGIT_WIDTH = 16;

const int SCORE_HEIGHT = 24;
const int SCORE_WIDTH = 108;

const int ATTEMPTS_HEIGHT = 30;
const int ATTEMPTS_WIDTH = 174;

const logic [10:0] PADDING = 5;

const logic [10:0] SCORE_H_X = SCORE_OFFSET_X + SCORE_WIDTH + PADDING;
const logic [10:0] SCORE_L_X = SCORE_OFFSET_X + SCORE_WIDTH + DIGIT_WIDTH + PADDING;
const logic [10:0] ATTEMPTS_H_X = ATTEMPTS_OFFSET_X + ATTEMPTS_WIDTH + PADDING;
const logic [10:0] ATTEMPTS_L_X = ATTEMPTS_OFFSET_X + ATTEMPTS_WIDTH + DIGIT_WIDTH + PADDING;

const logic [7:0] TRANSPARENT_ENCODING = 8'hff;
const logic [7:0] BLACK_ENCODING = 8'h00;
const logic [7:0] BLUE_ENCODING = 8'b00000011;
const logic [7:0] RED_ENCODING = 8'b11100000;


logic [10:0] offsetY;
logic [7:0] background;

always_ff @(posedge clk) begin
	RGBoutStat <= background;
	if(SCORE_OFFSET_X <= pixelX && pixelX < SCORE_OFFSET_X + SCORE_WIDTH && offsetY <= pixelY && pixelY < offsetY + SCORE_HEIGHT) begin
		RGBoutStat <= (SCORE_BITMAP[pixelY - offsetY][pixelX - SCORE_OFFSET_X]) ? BLUE_ENCODING : background;
	end
	else if(ATTEMPTS_OFFSET_X <= pixelX && pixelX < ATTEMPTS_OFFSET_X + ATTEMPTS_WIDTH && offsetY <= pixelY && pixelY < offsetY + ATTEMPTS_HEIGHT) begin
		RGBoutStat <= (ATTEMPTS_BITMAP[pixelY - offsetY][pixelX - ATTEMPTS_OFFSET_X]) ? RED_ENCODING : background;
	end
	
	else if (offsetY <= pixelY && pixelY < offsetY + DIGIT_HEIGHT) begin
		if(SCORE_H_X <= pixelX && pixelX < SCORE_H_X + DIGIT_WIDTH) begin
			RGBoutStat <= (DIGIT_BITMAP[score[7:4]][pixelY - offsetY][pixelX - SCORE_H_X]) ? BLUE_ENCODING : background;
		end
		else if(SCORE_L_X <= pixelX && pixelX < SCORE_L_X + DIGIT_WIDTH) begin
			RGBoutStat <= (DIGIT_BITMAP[score[3:0]][pixelY - offsetY][pixelX - SCORE_L_X]) ? BLUE_ENCODING : background;
		end
		else if(ATTEMPTS_H_X <= pixelX && pixelX < ATTEMPTS_H_X + DIGIT_WIDTH) begin
			RGBoutStat <= (DIGIT_BITMAP[attempts[7:4]][pixelY - offsetY][pixelX - ATTEMPTS_H_X]) ? RED_ENCODING : background;
		end
		else if(ATTEMPTS_L_X <= pixelX && pixelX < ATTEMPTS_L_X + DIGIT_WIDTH) begin
			RGBoutStat <= (DIGIT_BITMAP[attempts[3:0]][pixelY - offsetY][pixelX - ATTEMPTS_L_X]) ? RED_ENCODING : background;
		end
	end
	
end

always_comb begin
	if(gameFinished) begin
		offsetY = MIDDLE_OFFSET_Y;
		background = BLACK_ENCODING;
	end
	
	else begin
		offsetY = DOWN_OFFSET;
		background = TRANSPARENT_ENCODING;
	end
end

assign drawingRequestStat = (RGBoutStat != TRANSPARENT_ENCODING) ? 1'b1 : 1'b0;

logic[0:23][0:107] SCORE_BITMAP = {
	108'b000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	108'b000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	108'b001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	108'b011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	108'b011111110000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	108'b111111000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	108'b111111000000000001100000000001111111000000000001111111100000000001111100001110000000011111111000000000011111,
	108'b111111000000000000000000001111111111111000000111111111111000000001111100111110000001111111111110000000111111,
	108'b111111110000000000000000011111111111111000001111111111111100000001111111111110000011111111111111000000111111,
	108'b111111111111100000000000111111111111111000011111111111111110000001111111111110000111111111111111100000111111,
	108'b011111111111111100000001111111100001111000111111100001111111000001111111111110001111111000011111100000111111,
	108'b011111111111111110000001111110000000011000111111000000111111000001111110000000001111110000001111110000011111,
	108'b001111111111111111000001111110000000000000111111000000111111000001111100000000001111100000001111110000000000,
	108'b000011111111111111100001111100000000000001111110000000011111100001111100000000011111111111111111110000000000,
	108'b000000001111111111100011111100000000000001111110000000011111100001111100000000011111111111111111110000000000,
	108'b000000000000111111110011111100000000000001111110000000011111100001111100000000011111111111111111110000000000,
	108'b000000000000011111110011111100000000000001111110000000011111000001111100000000011111100000000000000000000000,
	108'b100000000000011111100001111110000000000000111111000000111111000001111100000000001111100000000000000000000000,
	108'b111000000000011111100001111110000000011000111111000000111111000001111100000000001111110000000000110000011111,
	108'b111111000000111111100001111111100000111000111111100001111111000001111100000000001111111100000011110000111111,
	108'b111111111111111111000000111111111111111000011111111111111110000001111100000000000111111111111111110000111111,
	108'b111111111111111110000000011111111111111000001111111111111100000001111100000000000011111111111111110000111111,
	108'b111111111111111100000000001111111111111000000111111111111000000001111100000000000001111111111111100000111111,
	108'b000011111111100000000000000001111111000000000001111111100000000001111100000000000000001111111110000000011111};
	
	logic[0:30][0:173] ATTEMPTS_BITMAP = {
	174'b000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
	174'b000000011111111000000000000111111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000,
	174'b000000011111111100000000000111111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000,
	174'b000000011111111100000000000111111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000,
	174'b000000111111111100000000000111111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000,
	174'b000000111111111110000000000111111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000,
	174'b000000111111111110000000011111111111110011111111111110000000001111111000000000111110001111100000001111100000000011111000111111000000111111111111100000001111111110000000011111,
	174'b000001111110111111000000011111111111110011111111111110000001111111111110000000111110011111111000111111111000000011111111111111100000111111111111100000111111111111100000111111,
	174'b000001111110111111000000011111111111110011111111111110000011111111111111000000111111111111111101111111111000000011111111111111110000111111111111100001111111111111100000111111,
	174'b000001111100111111000000011111111111110011111111111110000111111111111111100000111111111111111111111111111100000011111111111111111000111111111111100011111111111111100000111111,
	174'b000011111100011111100000000111111000000000111111000000001111111000011111100000111111111111111111111111111100000011111100001111111000001111110000000011111100000111100000111111,
	174'b000011111100011111100000000111111000000000111111000000001111110000001111110000111111000011111111000011111100000011111000000111111100001111110000000011111000000000100000011111,
	174'b000111111000011111100000000111111000000000111111000000001111100000001111110000111110000001111110000011111100000011111000000011111100001111110000000011111110000000000000000000,
	174'b000111111000001111110000000111111000000000111111000000011111111111111111110000111110000001111110000001111100000011111000000011111100001111110000000011111111111100000000000000,
	174'b000111111000001111110000000111111000000000111111000000011111111111111111110000111110000001111110000001111100000011111000000011111100001111110000000011111111111111000000000000,
	174'b001111111111111111110000000111111000000000111111000000011111111111111111110000111110000001111110000001111100000011111000000011111100001111110000000001111111111111100000000000,
	174'b001111111111111111111000000111111000000000111111000000011111100000000000000000111110000001111110000001111100000011111000000011111100001111110000000000011111111111110000000000,
	174'b001111111111111111111000000111111000000000111111000000001111100000000000000000111110000001111110000001111100000011111000000011111100001111110000000000000000111111110000000000,
	174'b011111111111111111111100000111111000000000111111000000001111110000000000110000111110000001111110000001111100000011111000000111111000001111110000000110000000001111110000011111,
	174'b011111100000000011111100000111111000010000111111000010001111111100000011110000111110000001111110000001111100000011111100001111111000001111110000100111110000001111110000111111,
	174'b011111100000000011111100000111111111110000111111111110000111111111111111110000111110000001111110000001111100000011111111111111110000001111111111100111111111111111100000111111,
	174'b111111000000000011111110000011111111110000011111111110000011111111111111110000111110000001111110000001111100000011111111111111110000000111111111100111111111111111100000111111,
	174'b111111000000000001111110000011111111110000011111111110000001111111111111100000111110000001111110000001111100000011111111111111000000000111111111100011111111111110000000111111,
	174'b111111000000000001111110000000111111100000000111111100000000001111111110000000111110000001111110000001111100000011111001111110000000000001111111000000111111111000000000011111,
	174'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000,
	174'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000,
	174'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000,
	174'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000,
	174'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000,
	174'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000};

logic [0:15] [0:31] [0:15] DIGIT_BITMAP = {
{16'b	0000001111100000,
16'b	0000111111111000,
16'b	0000111111111000,
16'b	0001111111111100,
16'b	0011111001111100,
16'b	0011100000111110,
16'b	0111100000011110,
16'b	0111100000011110,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000011110,
16'b	1111100000011110,
16'b	0111110000111110,
16'b	0111110000111100,
16'b	0011111001111100,
16'b	0011111111111000,
16'b	0001111111111000,
16'b	0000111111110000,
16'b	0000011111000000},

{16'b	0000000011100000,
16'b	0000000111100000,
16'b	0000011111100000,
16'b	0000111111100000,
16'b	0001111111100000,
16'b	0011111111100000,
16'b	0111111011100000,
16'b	0111100011100000,
16'b	0111000011100000,
16'b	0010000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111111},

{16'b	0000111111100000,
16'b	0001111111110000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000011111100,
16'b	1110000001111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000001111100,
16'b	0000000001111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011110000,
16'b	0000000011100000,
16'b	0000000111000000,
16'b	0000001111000000,
16'b	0000011110000000,
16'b	0000111100000000,
16'b	0001111100000000,
16'b	0001111100000000,
16'b	0011111000000000,
16'b	0111110000000001,
16'b	1111100000000011,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111},

{16'b	0000111111100000,
16'b	0001111111111000,
16'b	0111111111111000,
16'b	1111111111111000,
16'b	1111110011111100,
16'b	1111000001111100,
16'b	1110000001111100,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0001111111110000,
16'b	0001111111000000,
16'b	0001111111111000,
16'b	0001111111111000,
16'b	0000000011111100,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000111111,
16'b	1110000001111110,
16'b	1111100011111110,
16'b	1111111111111100,
16'b	1111111111111000,
16'b	0111111111111000,
16'b	0001111111000000},

{16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000111111000,
16'b	0000001111111000,
16'b	0000001101111000,
16'b	0000011101111000,
16'b	0000011101111000,
16'b	0000111101111000,
16'b	0001111101111000,
16'b	0001111101111000,
16'b	0001111001111000,
16'b	0011111001111000,
16'b	0011110001111000,
16'b	0111100001111000,
16'b	0111100001111000,
16'b	1111000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1110000001111000,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000001111000,
16'b	0000000011111100},

{16'b	0111111111111111,
16'b	0111111111111111,
16'b	0111111111111110,
16'b	0111111111111100,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	0111111111100000,
16'b	0111111111111000,
16'b	0111111111111000,
16'b	0111111111111100,
16'b	0010000011111110,
16'b	0000000001111110,
16'b	0000000000111111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000011111,
16'b	0000000000011111,
16'b	1000000000111110,
16'b	1100000001111110,
16'b	1111100011111100,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	0001111111000000},

{16'b	0000000111111100,
16'b	0000011111111110,
16'b	0000111111111110,
16'b	0001111111111111,
16'b	0001111100001111,
16'b	0011111100000001,
16'b	0011111000000000,
16'b	0111110000000000,
16'b	0111100000000000,
16'b	1111100000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111001111111000,
16'b	1111111111111100,
16'b	1111111111111110,
16'b	1111111111111111,
16'b	1111111101111111,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111000000000111,
16'b	1111100000001111,
16'b	1111100000001111,
16'b	0111110000011111,
16'b	0111111101111110,
16'b	0011111111111110,
16'b	0001111111111100,
16'b	0001111111111000,
16'b	0000011111100000},

{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1100000000001111,
16'b	1000000000011111,
16'b	0000000000011111,
16'b	0000000000011110,
16'b	0000000000111110,
16'b	0000000000111100,
16'b	0000000001111100,
16'b	0000000001111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011111000,
16'b	0000000011110000,
16'b	0000000011110000,
16'b	0000000011100000,
16'b	0000000011100000,
16'b	0000000111100000,
16'b	0000000111100000,
16'b	0000001111000000,
16'b	0000001111000000,
16'b	0000011110000000,
16'b	0000011110000000,
16'b	0000111110000000,
16'b	0000111100000000,
16'b	0000111100000000,
16'b	0001111100000000,
16'b	0001111100000000,
16'b	0001111100000000},

{16'b	0000111111110000,
16'b	0001111111111000,
16'b	0011111111111100,
16'b	0111111111111110,
16'b	0111111011111110,
16'b	1111100000111111,
16'b	1111100000011111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111000000001111,
16'b	1111100000011110,
16'b	0111110000111110,
16'b	0111111001111100,
16'b	0011111111111000,
16'b	0001111111111000,
16'b	0000111111100000,
16'b	0000111111110000,
16'b	0001111111111000,
16'b	0011111111111100,
16'b	0111111001111110,
16'b	1111100000111111,
16'b	1111000000001111,
16'b	1110000000001111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1111000000001111,
16'b	1111100000011111,
16'b	1111111001111111,
16'b	1111111111111110,
16'b	0111111111111110,
16'b	0011111111111000,
16'b	0001111111110000},
	
{16'b	0000111111100000,
16'b	0001111111111000,
16'b	0011111111111000,
16'b	0111111111111100,
16'b	1111111011111100,
16'b	1111100000111110,
16'b	1111000000011110,
16'b	1111000000011111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1110000000001111,
16'b	1111000000001111,
16'b	1111100000011111,
16'b	1111111011111111,
16'b	1111111111111111,
16'b	0111111111111111,
16'b	0011111111111111,
16'b	0001111111001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000001111,
16'b	0000000000011110,
16'b	0000000000011110,
16'b	0000000000111110,
16'b	0000000001111100,
16'b	1000000011111100,
16'b	1111000011111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	1111111111100000,
16'b	0011111100000000},

{16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000011111100000,
16'b	0000111111110000,
16'b	0000110000111000,
16'b	0000110000111000,
16'b	0000110000111000,
16'b	0001110000111100,
16'b	0001100000011100,
16'b	0011100000011100,
16'b	0011000000001100,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	0111000000001110,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1110000000000111,
16'b	1111000000001111},

{16'b	1111111111110000,
16'b	1111111111111000,
16'b	1111111111111100,
16'b	1111111111111110,
16'b	0111000011111110,
16'b	0111000000111111,
16'b	0111000000011111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000011110,
16'b	0111000000111110,
16'b	0111000001111100,
16'b	0111111111111000,
16'b	0111111111111000,
16'b	0111111111100000,
16'b	0111111111110000,
16'b	0111111111111000,
16'b	0111111111111100,
16'b	0111000001111110,
16'b	0111000000111111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000000111,
16'b	0111000000000111,
16'b	0111000000001111,
16'b	0111000000011111,
16'b	0111000001111111,
16'b	1111111111111110,
16'b	1111111111111110,
16'b	1111111111111000,
16'b	1111111111110000},

{16'b	0000001111111000,
16'b	0000111111111100,
16'b	0000111111111110,
16'b	0001111111111111,
16'b	0011111001000011,
16'b	0011100000000001,
16'b	0111100000000000,
16'b	0111100000000000,
16'b	1111100000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111100000000000,
16'b	0111110000000000,
16'b	0111110000000001,
16'b	0011111001000011,
16'b	0011111111111111,
16'b	0001111111111110,
16'b	0000111111111100,
16'b	0000011111111000},

{16'b	1111111111100000,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111111100,
16'b	0111000001111100,
16'b	0111000000111110,
16'b	0111000000011110,
16'b	0111000000011110,
16'b	0111000000011111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000001111,
16'b	0111000000011110,
16'b	0111000000011110,
16'b	0111000000111110,
16'b	0111000000111100,
16'b	0111000001111100,
16'b	1111111111111000,
16'b	1111111111111000,
16'b	1111111111110000,
16'b	1111111111000000},

{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000011,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000001,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000001,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000001000011,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111},

{16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000011,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000001,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111111111111111,
16'b	1111000000000001,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000,
16'b	1111000000000000}};

endmodule
