module holes (
					input logic clk,
					input logic resetN,
					input logic signed [10:0] pixelX,
					input logic signed [10:0] pixelY,

					output logic drawingRequestHoles,
					output logic [7:0] RGBoutHoles
);


endmodule
